
interface bus_if (input pclk, input presetn);
	//declare interface signals
  
endinterface
