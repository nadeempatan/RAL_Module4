// Declare a sequence_item for the APB transaction
class cretae bus_pkt class extended from uvm_sequence_item


//function new	
endclass
/////////////////////
