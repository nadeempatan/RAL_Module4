
// Monitors the APB interface for any activity and reports out
// through an analysis port
class create monitor clas extended from uvm_monitor
//factroy registration
//

//declare analysis port and virtual interface

//function new
//
//
//
//

//run phase
  virtual task run_phase (uvm_phase phase);





  endtask
endclass
