
// Register environment class puts together the model,adapter and predictor
class create ral_env  extended from uvm_env
 `uvm_component_utils (reg_env)
 //function new


 //register model handle
 //adapter 
 //predictor handle
 
 //buildphase

 //create instance for model adapter and predictor
 //
 //
 
 //build model
 //
 
 //lock model
 //
 /


  //connect phase

//connect predictor to map
//

//connect predictor to adapter
//

// connect predictor to mointor analysis port


endclass
/////////
