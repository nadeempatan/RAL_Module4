class //create sequencer class seqcr extended from uvm sequencer
// factory registration
//
//
//

//function new
  
 

//build phase
endclass
