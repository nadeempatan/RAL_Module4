//include all the files inside pacakage 
//
//
//

/*`include "transaction.sv"
`include "sequencer.sv"
`include "monitor.sv"
`include "driver.sv"
`include "agent.sv"
`include "base_seq.sv"
`include "reg_model.sv"
`include "reg2apb_adaptor.sv"
`include "ral_env.sv"
`include "env.sv"
`include "base_test.sv"

*/
