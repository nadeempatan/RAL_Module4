// Drives a given apb transaction packet to the APB interface
class create driver clas extended from uvm driver
 // factory registration
 

 //tarnsaction and virtual interface handle
 //
 //
 
 //function new
 //
 //
 //
 //
 
 //build pahse
 //
 //
 //
 //
 
 //run pahse
   virtual task run_phase (uvm_phase phase);



 endtask
endclass
