// The agent puts together the driver, sequencer and monitor 
class //create agent class extended from uvm_agent;
 // registration 
 //
 
// handle of driver sequencer and monitor

 //function new
 //

 //build phase


 // create an instance for driver ,sequencer and moitor

 //connect phase
endclass
