class//create env class extended from uvm_env class


//factory registration
 

 // agent handle
 // reg env handle
 //
 
 //function new


// build phase 

 //cretae an instance of agent and reg env
 //
 //
 //
 
 

//connect phase
 // Connect analysis port of monitor with predictor, assign agent to register env
 // and set default map of the register env
//inside connect function
 //connect analysis port of monitor with predictor
 //set default map of the reg_env

endclass
