
class //create testclass  extended from uvm_test
 // factroy registration 
 

//env handle 
//
//
//

//function new


//build phase
// Build the testbench environment 


 //run phase
 //start seq
endclass
