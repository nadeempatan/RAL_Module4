class //create seq extends uvm_sequence
//factory registration 
//
//
//

//function new
  
//task body
  task body();

   endtask
endclass
